* File: 4_bit_accumulator.pex.netlist
* Created: Mon Nov  9 17:56:30 2020
* Program "Calibre xRC"
* Version "v2011.3_29.20"
* 

* Transistor models.
.include '$PDK_DIR/ncsu_basekit/models/hspice/hspice_nom.include'

* Analysis commands
.param vdd_val = 1.1
.param clk_period = 100
.param rise_fall_time = 0.10 * clk_period

Vsupply vdd 0 vdd_val
Vgnd gnd 0 0

* Digital vector file for input from same directory
.vec '4bit_input.vec'

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    POST

.include "4_bit_accumulator.pex.netlist.pex"

.subckt 4_bit_accumulator  GND PHI RST VDD CIN COUT A0 SOUT0 A1 SOUT1 A2 SOUT2
+ A3 SOUT3
* 
* SOUT3	SOUT3
* A3	A3
* SOUT2	SOUT2
* A2	A2
* SOUT1	SOUT1
* A1	A1
* SOUT0	SOUT0
* A0	A0
* COUT	COUT
* CIN	CIN
* VDD	VDD
* RST	RST
* PHI	PHI
* GND	GND
mXI0/XI0/XI0/MM0 N_NET5_XI0/XI0/XI0/MM0_d N_XI0/XI0/NET20_XI0/XI0/XI0/MM0_g
+ N_XI0/XI0/XI0/NET15_XI0/XI0/XI0/MM0_s N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI0/XI0/XI0/MM3 N_XI0/XI0/XI0/NET15_XI0/XI0/XI0/MM3_d
+ N_XI0/XI0/NET19_XI0/XI0/XI0/MM3_g N_GND_XI0/XI0/XI0/MM3_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI0/XI0/MM2 N_XI0/XI0/XI0/NET15_XI0/XI0/XI0/MM3_d
+ N_XI0/XI0/NET18_XI0/XI0/XI0/MM2_g N_GND_XI0/XI0/XI0/MM2_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI1/MM0 N_XI0/NET20_XI0/XI1/MM0_d N_XI0/NET21_XI0/XI1/MM0_g
+ N_VDD_XI0/XI1/MM0_s N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI0/XI1/MM1 N_XI0/NET20_XI0/XI1/MM0_d N_RST_XI0/XI1/MM1_g N_VDD_XI0/XI1/MM1_s
+ N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI0/XI0/MM5 N_NET5_XI0/XI0/XI0/MM5_d N_XI0/XI0/NET20_XI0/XI0/XI0/MM5_g
+ N_XI0/XI0/XI0/NET17_XI0/XI0/XI0/MM5_s N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08
+ W=3.6e-07 AD=3.78e-14 AS=3.78e-14 PD=9.3e-07 PS=9.3e-07
mXI0/XI0/XI0/MM8 N_XI0/XI0/XI0/NET17_XI0/XI0/XI0/MM8_d
+ N_XI0/XI0/NET19_XI0/XI0/XI0/MM8_g N_VDD_XI0/XI0/XI0/MM8_s
+ N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI0/XI0/XI0/MM7 N_XI0/XI0/XI0/NET17_XI0/XI0/XI0/MM8_d
+ N_XI0/XI0/NET18_XI0/XI0/XI0/MM7_g N_VDD_XI0/XI0/XI0/MM7_s
+ N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI0/XI0/XI1/MM6 N_XI0/XI0/XI1/NET26_XI0/XI0/XI1/MM6_d N_A0_XI0/XI0/XI1/MM6_g
+ N_VDD_XI0/XI0/XI1/MM6_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07
+ AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI0/XI0/XI1/MM7 N_XI0/XI0/XI1/NET32_XI0/XI0/XI1/MM7_d
+ N_XI0/XI0/NET18_XI0/XI0/XI1/MM7_g N_VDD_XI0/XI0/XI1/MM7_s
+ N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=5.67e-14
+ PD=1.29e-06 PS=1.29e-06
mXI0/XI0/XI1/MM0 N_XI0/NET21_XI0/XI0/XI1/MM0_d N_XI0/XI0/NET20_XI0/XI0/XI1/MM0_g
+ N_XI0/XI0/XI1/NET25_XI0/XI0/XI1/MM0_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI0/XI0/XI1/MM1 N_XI0/NET21_XI0/XI0/XI1/MM1_d N_CIN_XI0/XI0/XI1/MM1_g
+ N_XI0/XI0/XI1/NET31_XI0/XI0/XI1/MM1_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI0/XI0/XI1/MM14 N_XI0/XI0/XI1/NET22_XI0/XI0/XI1/MM14_d N_A0_XI0/XI0/XI1/MM14_g
+ N_GND_XI0/XI0/XI1/MM14_s N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07
+ AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI0/XI0/XI1/MM15 N_XI0/XI0/XI1/NET28_XI0/XI0/XI1/MM15_d
+ N_XI0/XI0/NET18_XI0/XI0/XI1/MM15_g N_GND_XI0/XI0/XI1/MM15_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14
+ PD=7.5e-07 PS=7.5e-07
mXI0/XI0/XI1/MM8 N_XI0/NET21_XI0/XI0/XI1/MM8_d N_XI0/XI0/NET20_XI0/XI0/XI1/MM8_g
+ N_XI0/XI0/XI1/NET23_XI0/XI0/XI1/MM8_s N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI0/XI0/XI1/MM9 N_XI0/NET21_XI0/XI0/XI1/MM9_d N_CIN_XI0/XI0/XI1/MM9_g
+ N_XI0/XI0/XI1/NET29_XI0/XI0/XI1/MM9_s N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI0/XI0/XI3/MM0 N_XI0/XI0/NET18_XI0/XI0/XI3/MM0_d N_A0_XI0/XI0/XI3/MM0_g
+ N_GND_XI0/XI0/XI3/MM0_s N_GND_XI0/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI0/XI2/XI4/MM0 N_XI0/XI2/NET22_XI0/XI2/XI4/MM0_d N_PHI_XI0/XI2/XI4/MM0_g
+ N_GND_XI0/XI2/XI4/MM0_s N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI0/XI0/XI4/MM0 N_XI0/XI0/NET19_XI0/XI0/XI4/MM0_d N_SOUT0_XI0/XI0/XI4/MM0_g
+ N_GND_XI0/XI0/XI4/MM0_s N_GND_XI0/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI0/XI2/XI3/MM0 N_SOUT0_XI0/XI2/XI3/MM0_d N_XI0/XI2/NET17_XI0/XI2/XI3/MM0_g
+ N_GND_XI0/XI2/XI3/MM0_s N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI0/XI0/XI2/MM0 N_XI0/XI0/NET20_XI0/XI0/XI2/MM0_d N_CIN_XI0/XI0/XI2/MM0_g
+ N_GND_XI0/XI0/XI2/MM0_s N_GND_XI0/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI0/XI0/XI3/MM1 N_XI0/XI0/NET18_XI0/XI0/XI3/MM1_d N_A0_XI0/XI0/XI3/MM1_g
+ N_VDD_XI0/XI0/XI3/MM1_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI0/XI2/XI4/MM1 N_XI0/XI2/NET22_XI0/XI2/XI4/MM1_d N_PHI_XI0/XI2/XI4/MM1_g
+ N_VDD_XI0/XI2/XI4/MM1_s N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI0/XI0/XI4/MM1 N_XI0/XI0/NET19_XI0/XI0/XI4/MM1_d N_SOUT0_XI0/XI0/XI4/MM1_g
+ N_VDD_XI0/XI0/XI4/MM1_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI0/XI2/XI3/MM1 N_SOUT0_XI0/XI2/XI3/MM1_d N_XI0/XI2/NET17_XI0/XI2/XI3/MM1_g
+ N_VDD_XI0/XI2/XI3/MM1_s N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI0/XI0/XI2/MM1 N_XI0/XI0/NET20_XI0/XI0/XI2/MM1_d N_CIN_XI0/XI0/XI2/MM1_g
+ N_VDD_XI0/XI0/XI2/MM1_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI0/XI0/XI1/MM3 N_XI0/XI0/XI1/NET25_XI0/XI0/XI1/MM3_d
+ N_XI0/XI0/NET19_XI0/XI0/XI1/MM3_g N_XI0/XI0/XI1/NET32_XI0/XI0/XI1/MM3_s
+ N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI0/XI0/XI1/MM2 N_XI0/XI0/XI1/NET25_XI0/XI0/XI1/MM3_d N_SOUT0_XI0/XI0/XI1/MM2_g
+ N_XI0/XI0/XI1/NET26_XI0/XI0/XI1/MM2_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI0/XI0/XI1/MM5 N_XI0/XI0/XI1/NET31_XI0/XI0/XI1/MM5_d N_SOUT0_XI0/XI0/XI1/MM5_g
+ N_XI0/XI0/XI1/NET32_XI0/XI0/XI1/MM5_s N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI0/XI0/XI1/MM4 N_XI0/XI0/XI1/NET31_XI0/XI0/XI1/MM5_d
+ N_XI0/XI0/NET19_XI0/XI0/XI1/MM4_g N_XI0/XI0/XI1/NET26_XI0/XI0/XI1/MM4_s
+ N_VDD_XI0/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI0/XI0/XI1/MM11 N_XI0/XI0/XI1/NET23_XI0/XI0/XI1/MM11_d
+ N_XI0/XI0/NET19_XI0/XI0/XI1/MM11_g N_XI0/XI0/XI1/NET28_XI0/XI0/XI1/MM11_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI0/XI0/XI1/MM10 N_XI0/XI0/XI1/NET23_XI0/XI0/XI1/MM11_d
+ N_SOUT0_XI0/XI0/XI1/MM10_g N_XI0/XI0/XI1/NET22_XI0/XI0/XI1/MM10_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI0/XI0/XI1/MM13 N_XI0/XI0/XI1/NET29_XI0/XI0/XI1/MM13_d
+ N_SOUT0_XI0/XI0/XI1/MM13_g N_XI0/XI0/XI1/NET28_XI0/XI0/XI1/MM13_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI0/XI0/XI1/MM12 N_XI0/XI0/XI1/NET29_XI0/XI0/XI1/MM13_d
+ N_XI0/XI0/NET19_XI0/XI0/XI1/MM12_g N_XI0/XI0/XI1/NET22_XI0/XI0/XI1/MM12_s
+ N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI0/XI0/XI0/MM9 XI0/XI0/XI0/NET30 N_XI0/XI0/NET19_XI0/XI0/XI0/MM9_g
+ N_VDD_XI0/XI0/XI0/MM9_s N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=5.04e-14 AS=3.78e-14 PD=1e-06 PS=9.3e-07
mXI0/XI0/XI0/MM6 N_NET5_XI0/XI0/XI0/MM6_d N_XI0/XI0/NET18_XI0/XI0/XI0/MM6_g
+ XI0/XI0/XI0/NET30 N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=3.78e-14 AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI0/XI2/MM7 XI0/XI2/NET29 N_XI0/NET20_XI0/XI2/MM7_g N_VDD_XI0/XI2/MM7_s
+ N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI0/XI2/MM6 N_XI0/XI2/NET15_XI0/XI2/MM6_d N_PHI_XI0/XI2/MM6_g XI0/XI2/NET29
+ N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
mXI0/XI2/MM5 XI0/XI2/NET28 N_XI0/XI2/NET15_XI0/XI2/MM5_g N_VDD_XI0/XI2/MM5_s
+ N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI0/XI2/MM4 N_XI0/XI2/NET17_XI0/XI2/MM4_d N_XI0/XI2/NET22_XI0/XI2/MM4_g
+ XI0/XI2/NET28 N_VDD_XI0/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14
+ AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI0/XI1/MM3 XI0/XI1/NET15 N_XI0/NET21_XI0/XI1/MM3_g N_GND_XI0/XI1/MM3_s
+ N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI1/MM2 N_XI0/NET20_XI0/XI1/MM2_d N_RST_XI0/XI1/MM2_g XI0/XI1/NET15
+ N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI0/XI0/XI0/MM4 XI0/XI0/XI0/NET29 N_XI0/XI0/NET19_XI0/XI0/XI0/MM4_g
+ N_GND_XI0/XI0/XI0/MM4_s N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI0/XI0/XI0/MM1 N_NET5_XI0/XI0/XI0/MM1_d N_XI0/XI0/NET18_XI0/XI0/XI0/MM1_g
+ XI0/XI0/XI0/NET29 N_GND_XI0/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI0/XI2/MM1 XI0/XI2/NET26 N_XI0/NET20_XI0/XI2/MM1_g N_GND_XI0/XI2/MM1_s
+ N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI2/MM8 N_XI0/XI2/NET15_XI0/XI2/MM8_d N_XI0/XI2/NET22_XI0/XI2/MM8_g
+ XI0/XI2/NET26 N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14
+ AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI0/XI2/MM2 XI0/XI2/NET023 N_XI0/XI2/NET15_XI0/XI2/MM2_g N_GND_XI0/XI2/MM2_s
+ N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI0/XI2/MM0 N_XI0/XI2/NET17_XI0/XI2/MM0_d N_PHI_XI0/XI2/MM0_g XI0/XI2/NET023
+ N_GND_XI0/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI0/XI0/MM0 N_NET4_XI1/XI0/XI0/MM0_d N_XI1/XI0/NET20_XI1/XI0/XI0/MM0_g
+ N_XI1/XI0/XI0/NET15_XI1/XI0/XI0/MM0_s N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI1/XI0/XI0/MM3 N_XI1/XI0/XI0/NET15_XI1/XI0/XI0/MM3_d
+ N_XI1/XI0/NET19_XI1/XI0/XI0/MM3_g N_GND_XI1/XI0/XI0/MM3_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI0/XI0/MM2 N_XI1/XI0/XI0/NET15_XI1/XI0/XI0/MM3_d
+ N_XI1/XI0/NET18_XI1/XI0/XI0/MM2_g N_GND_XI1/XI0/XI0/MM2_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI1/MM0 N_XI1/NET20_XI1/XI1/MM0_d N_XI1/NET21_XI1/XI1/MM0_g
+ N_VDD_XI1/XI1/MM0_s N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI1/XI1/MM1 N_XI1/NET20_XI1/XI1/MM0_d N_RST_XI1/XI1/MM1_g N_VDD_XI1/XI1/MM1_s
+ N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI0/XI0/MM5 N_NET4_XI1/XI0/XI0/MM5_d N_XI1/XI0/NET20_XI1/XI0/XI0/MM5_g
+ N_XI1/XI0/XI0/NET17_XI1/XI0/XI0/MM5_s N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08
+ W=3.6e-07 AD=3.78e-14 AS=3.78e-14 PD=9.3e-07 PS=9.3e-07
mXI1/XI0/XI0/MM8 N_XI1/XI0/XI0/NET17_XI1/XI0/XI0/MM8_d
+ N_XI1/XI0/NET19_XI1/XI0/XI0/MM8_g N_VDD_XI1/XI0/XI0/MM8_s
+ N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI1/XI0/XI0/MM7 N_XI1/XI0/XI0/NET17_XI1/XI0/XI0/MM8_d
+ N_XI1/XI0/NET18_XI1/XI0/XI0/MM7_g N_VDD_XI1/XI0/XI0/MM7_s
+ N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI1/XI0/XI1/MM6 N_XI1/XI0/XI1/NET26_XI1/XI0/XI1/MM6_d N_A1_XI1/XI0/XI1/MM6_g
+ N_VDD_XI1/XI0/XI1/MM6_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07
+ AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI1/XI0/XI1/MM7 N_XI1/XI0/XI1/NET32_XI1/XI0/XI1/MM7_d
+ N_XI1/XI0/NET18_XI1/XI0/XI1/MM7_g N_VDD_XI1/XI0/XI1/MM7_s
+ N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=5.67e-14
+ PD=1.29e-06 PS=1.29e-06
mXI1/XI0/XI1/MM0 N_XI1/NET21_XI1/XI0/XI1/MM0_d N_XI1/XI0/NET20_XI1/XI0/XI1/MM0_g
+ N_XI1/XI0/XI1/NET25_XI1/XI0/XI1/MM0_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI1/XI0/XI1/MM1 N_XI1/NET21_XI1/XI0/XI1/MM1_d N_NET5_XI1/XI0/XI1/MM1_g
+ N_XI1/XI0/XI1/NET31_XI1/XI0/XI1/MM1_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI1/XI0/XI1/MM14 N_XI1/XI0/XI1/NET22_XI1/XI0/XI1/MM14_d N_A1_XI1/XI0/XI1/MM14_g
+ N_GND_XI1/XI0/XI1/MM14_s N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07
+ AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI1/XI0/XI1/MM15 N_XI1/XI0/XI1/NET28_XI1/XI0/XI1/MM15_d
+ N_XI1/XI0/NET18_XI1/XI0/XI1/MM15_g N_GND_XI1/XI0/XI1/MM15_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14
+ PD=7.5e-07 PS=7.5e-07
mXI1/XI0/XI1/MM8 N_XI1/NET21_XI1/XI0/XI1/MM8_d N_XI1/XI0/NET20_XI1/XI0/XI1/MM8_g
+ N_XI1/XI0/XI1/NET23_XI1/XI0/XI1/MM8_s N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI1/XI0/XI1/MM9 N_XI1/NET21_XI1/XI0/XI1/MM9_d N_NET5_XI1/XI0/XI1/MM9_g
+ N_XI1/XI0/XI1/NET29_XI1/XI0/XI1/MM9_s N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI1/XI0/XI3/MM0 N_XI1/XI0/NET18_XI1/XI0/XI3/MM0_d N_A1_XI1/XI0/XI3/MM0_g
+ N_GND_XI1/XI0/XI3/MM0_s N_GND_XI1/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI1/XI2/XI4/MM0 N_XI1/XI2/NET22_XI1/XI2/XI4/MM0_d N_PHI_XI1/XI2/XI4/MM0_g
+ N_GND_XI1/XI2/XI4/MM0_s N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI1/XI0/XI4/MM0 N_XI1/XI0/NET19_XI1/XI0/XI4/MM0_d N_SOUT1_XI1/XI0/XI4/MM0_g
+ N_GND_XI1/XI0/XI4/MM0_s N_GND_XI1/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI1/XI2/XI3/MM0 N_SOUT1_XI1/XI2/XI3/MM0_d N_XI1/XI2/NET17_XI1/XI2/XI3/MM0_g
+ N_GND_XI1/XI2/XI3/MM0_s N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI1/XI0/XI2/MM0 N_XI1/XI0/NET20_XI1/XI0/XI2/MM0_d N_NET5_XI1/XI0/XI2/MM0_g
+ N_GND_XI1/XI0/XI2/MM0_s N_GND_XI1/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI1/XI0/XI3/MM1 N_XI1/XI0/NET18_XI1/XI0/XI3/MM1_d N_A1_XI1/XI0/XI3/MM1_g
+ N_VDD_XI1/XI0/XI3/MM1_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI1/XI2/XI4/MM1 N_XI1/XI2/NET22_XI1/XI2/XI4/MM1_d N_PHI_XI1/XI2/XI4/MM1_g
+ N_VDD_XI1/XI2/XI4/MM1_s N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI1/XI0/XI4/MM1 N_XI1/XI0/NET19_XI1/XI0/XI4/MM1_d N_SOUT1_XI1/XI0/XI4/MM1_g
+ N_VDD_XI1/XI0/XI4/MM1_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI1/XI2/XI3/MM1 N_SOUT1_XI1/XI2/XI3/MM1_d N_XI1/XI2/NET17_XI1/XI2/XI3/MM1_g
+ N_VDD_XI1/XI2/XI3/MM1_s N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI1/XI0/XI2/MM1 N_XI1/XI0/NET20_XI1/XI0/XI2/MM1_d N_NET5_XI1/XI0/XI2/MM1_g
+ N_VDD_XI1/XI0/XI2/MM1_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI1/XI0/XI1/MM3 N_XI1/XI0/XI1/NET25_XI1/XI0/XI1/MM3_d
+ N_XI1/XI0/NET19_XI1/XI0/XI1/MM3_g N_XI1/XI0/XI1/NET32_XI1/XI0/XI1/MM3_s
+ N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI1/XI0/XI1/MM2 N_XI1/XI0/XI1/NET25_XI1/XI0/XI1/MM3_d N_SOUT1_XI1/XI0/XI1/MM2_g
+ N_XI1/XI0/XI1/NET26_XI1/XI0/XI1/MM2_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI1/XI0/XI1/MM5 N_XI1/XI0/XI1/NET31_XI1/XI0/XI1/MM5_d N_SOUT1_XI1/XI0/XI1/MM5_g
+ N_XI1/XI0/XI1/NET32_XI1/XI0/XI1/MM5_s N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI1/XI0/XI1/MM4 N_XI1/XI0/XI1/NET31_XI1/XI0/XI1/MM5_d
+ N_XI1/XI0/NET19_XI1/XI0/XI1/MM4_g N_XI1/XI0/XI1/NET26_XI1/XI0/XI1/MM4_s
+ N_VDD_XI1/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI1/XI0/XI1/MM11 N_XI1/XI0/XI1/NET23_XI1/XI0/XI1/MM11_d
+ N_XI1/XI0/NET19_XI1/XI0/XI1/MM11_g N_XI1/XI0/XI1/NET28_XI1/XI0/XI1/MM11_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI1/XI0/XI1/MM10 N_XI1/XI0/XI1/NET23_XI1/XI0/XI1/MM11_d
+ N_SOUT1_XI1/XI0/XI1/MM10_g N_XI1/XI0/XI1/NET22_XI1/XI0/XI1/MM10_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI1/XI0/XI1/MM13 N_XI1/XI0/XI1/NET29_XI1/XI0/XI1/MM13_d
+ N_SOUT1_XI1/XI0/XI1/MM13_g N_XI1/XI0/XI1/NET28_XI1/XI0/XI1/MM13_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI1/XI0/XI1/MM12 N_XI1/XI0/XI1/NET29_XI1/XI0/XI1/MM13_d
+ N_XI1/XI0/NET19_XI1/XI0/XI1/MM12_g N_XI1/XI0/XI1/NET22_XI1/XI0/XI1/MM12_s
+ N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI1/XI0/XI0/MM9 XI1/XI0/XI0/NET30 N_XI1/XI0/NET19_XI1/XI0/XI0/MM9_g
+ N_VDD_XI1/XI0/XI0/MM9_s N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=5.04e-14 AS=3.78e-14 PD=1e-06 PS=9.3e-07
mXI1/XI0/XI0/MM6 N_NET4_XI1/XI0/XI0/MM6_d N_XI1/XI0/NET18_XI1/XI0/XI0/MM6_g
+ XI1/XI0/XI0/NET30 N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=3.78e-14 AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI1/XI2/MM7 XI1/XI2/NET29 N_XI1/NET20_XI1/XI2/MM7_g N_VDD_XI1/XI2/MM7_s
+ N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI1/XI2/MM6 N_XI1/XI2/NET15_XI1/XI2/MM6_d N_PHI_XI1/XI2/MM6_g XI1/XI2/NET29
+ N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
mXI1/XI2/MM5 XI1/XI2/NET28 N_XI1/XI2/NET15_XI1/XI2/MM5_g N_VDD_XI1/XI2/MM5_s
+ N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI1/XI2/MM4 N_XI1/XI2/NET17_XI1/XI2/MM4_d N_XI1/XI2/NET22_XI1/XI2/MM4_g
+ XI1/XI2/NET28 N_VDD_XI1/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14
+ AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI1/XI1/MM3 XI1/XI1/NET15 N_XI1/NET21_XI1/XI1/MM3_g N_GND_XI1/XI1/MM3_s
+ N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI1/MM2 N_XI1/NET20_XI1/XI1/MM2_d N_RST_XI1/XI1/MM2_g XI1/XI1/NET15
+ N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI1/XI0/XI0/MM4 XI1/XI0/XI0/NET29 N_XI1/XI0/NET19_XI1/XI0/XI0/MM4_g
+ N_GND_XI1/XI0/XI0/MM4_s N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI1/XI0/XI0/MM1 N_NET4_XI1/XI0/XI0/MM1_d N_XI1/XI0/NET18_XI1/XI0/XI0/MM1_g
+ XI1/XI0/XI0/NET29 N_GND_XI1/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI1/XI2/MM1 XI1/XI2/NET26 N_XI1/NET20_XI1/XI2/MM1_g N_GND_XI1/XI2/MM1_s
+ N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI2/MM8 N_XI1/XI2/NET15_XI1/XI2/MM8_d N_XI1/XI2/NET22_XI1/XI2/MM8_g
+ XI1/XI2/NET26 N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14
+ AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI1/XI2/MM2 XI1/XI2/NET023 N_XI1/XI2/NET15_XI1/XI2/MM2_g N_GND_XI1/XI2/MM2_s
+ N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI1/XI2/MM0 N_XI1/XI2/NET17_XI1/XI2/MM0_d N_PHI_XI1/XI2/MM0_g XI1/XI2/NET023
+ N_GND_XI1/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI0/XI0/MM0 N_NET3_XI2/XI0/XI0/MM0_d N_XI2/XI0/NET20_XI2/XI0/XI0/MM0_g
+ N_XI2/XI0/XI0/NET15_XI2/XI0/XI0/MM0_s N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI2/XI0/XI0/MM3 N_XI2/XI0/XI0/NET15_XI2/XI0/XI0/MM3_d
+ N_XI2/XI0/NET19_XI2/XI0/XI0/MM3_g N_GND_XI2/XI0/XI0/MM3_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI0/XI0/MM2 N_XI2/XI0/XI0/NET15_XI2/XI0/XI0/MM3_d
+ N_XI2/XI0/NET18_XI2/XI0/XI0/MM2_g N_GND_XI2/XI0/XI0/MM2_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI1/MM0 N_XI2/NET20_XI2/XI1/MM0_d N_XI2/NET21_XI2/XI1/MM0_g
+ N_VDD_XI2/XI1/MM0_s N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI2/XI1/MM1 N_XI2/NET20_XI2/XI1/MM0_d N_RST_XI2/XI1/MM1_g N_VDD_XI2/XI1/MM1_s
+ N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI0/XI0/MM5 N_NET3_XI2/XI0/XI0/MM5_d N_XI2/XI0/NET20_XI2/XI0/XI0/MM5_g
+ N_XI2/XI0/XI0/NET17_XI2/XI0/XI0/MM5_s N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08
+ W=3.6e-07 AD=3.78e-14 AS=3.78e-14 PD=9.3e-07 PS=9.3e-07
mXI2/XI0/XI0/MM8 N_XI2/XI0/XI0/NET17_XI2/XI0/XI0/MM8_d
+ N_XI2/XI0/NET19_XI2/XI0/XI0/MM8_g N_VDD_XI2/XI0/XI0/MM8_s
+ N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI2/XI0/XI0/MM7 N_XI2/XI0/XI0/NET17_XI2/XI0/XI0/MM8_d
+ N_XI2/XI0/NET18_XI2/XI0/XI0/MM7_g N_VDD_XI2/XI0/XI0/MM7_s
+ N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI2/XI0/XI1/MM6 N_XI2/XI0/XI1/NET26_XI2/XI0/XI1/MM6_d N_A2_XI2/XI0/XI1/MM6_g
+ N_VDD_XI2/XI0/XI1/MM6_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07
+ AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI2/XI0/XI1/MM7 N_XI2/XI0/XI1/NET32_XI2/XI0/XI1/MM7_d
+ N_XI2/XI0/NET18_XI2/XI0/XI1/MM7_g N_VDD_XI2/XI0/XI1/MM7_s
+ N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=5.67e-14
+ PD=1.29e-06 PS=1.29e-06
mXI2/XI0/XI1/MM0 N_XI2/NET21_XI2/XI0/XI1/MM0_d N_XI2/XI0/NET20_XI2/XI0/XI1/MM0_g
+ N_XI2/XI0/XI1/NET25_XI2/XI0/XI1/MM0_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI2/XI0/XI1/MM1 N_XI2/NET21_XI2/XI0/XI1/MM1_d N_NET4_XI2/XI0/XI1/MM1_g
+ N_XI2/XI0/XI1/NET31_XI2/XI0/XI1/MM1_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI2/XI0/XI1/MM14 N_XI2/XI0/XI1/NET22_XI2/XI0/XI1/MM14_d N_A2_XI2/XI0/XI1/MM14_g
+ N_GND_XI2/XI0/XI1/MM14_s N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07
+ AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI2/XI0/XI1/MM15 N_XI2/XI0/XI1/NET28_XI2/XI0/XI1/MM15_d
+ N_XI2/XI0/NET18_XI2/XI0/XI1/MM15_g N_GND_XI2/XI0/XI1/MM15_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14
+ PD=7.5e-07 PS=7.5e-07
mXI2/XI0/XI1/MM8 N_XI2/NET21_XI2/XI0/XI1/MM8_d N_XI2/XI0/NET20_XI2/XI0/XI1/MM8_g
+ N_XI2/XI0/XI1/NET23_XI2/XI0/XI1/MM8_s N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI2/XI0/XI1/MM9 N_XI2/NET21_XI2/XI0/XI1/MM9_d N_NET4_XI2/XI0/XI1/MM9_g
+ N_XI2/XI0/XI1/NET29_XI2/XI0/XI1/MM9_s N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI2/XI0/XI3/MM0 N_XI2/XI0/NET18_XI2/XI0/XI3/MM0_d N_A2_XI2/XI0/XI3/MM0_g
+ N_GND_XI2/XI0/XI3/MM0_s N_GND_XI2/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI2/XI2/XI4/MM0 N_XI2/XI2/NET22_XI2/XI2/XI4/MM0_d N_PHI_XI2/XI2/XI4/MM0_g
+ N_GND_XI2/XI2/XI4/MM0_s N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI2/XI0/XI4/MM0 N_XI2/XI0/NET19_XI2/XI0/XI4/MM0_d N_SOUT2_XI2/XI0/XI4/MM0_g
+ N_GND_XI2/XI0/XI4/MM0_s N_GND_XI2/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI2/XI2/XI3/MM0 N_SOUT2_XI2/XI2/XI3/MM0_d N_XI2/XI2/NET17_XI2/XI2/XI3/MM0_g
+ N_GND_XI2/XI2/XI3/MM0_s N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI2/XI0/XI2/MM0 N_XI2/XI0/NET20_XI2/XI0/XI2/MM0_d N_NET4_XI2/XI0/XI2/MM0_g
+ N_GND_XI2/XI0/XI2/MM0_s N_GND_XI2/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI2/XI0/XI3/MM1 N_XI2/XI0/NET18_XI2/XI0/XI3/MM1_d N_A2_XI2/XI0/XI3/MM1_g
+ N_VDD_XI2/XI0/XI3/MM1_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI2/XI2/XI4/MM1 N_XI2/XI2/NET22_XI2/XI2/XI4/MM1_d N_PHI_XI2/XI2/XI4/MM1_g
+ N_VDD_XI2/XI2/XI4/MM1_s N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI2/XI0/XI4/MM1 N_XI2/XI0/NET19_XI2/XI0/XI4/MM1_d N_SOUT2_XI2/XI0/XI4/MM1_g
+ N_VDD_XI2/XI0/XI4/MM1_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI2/XI2/XI3/MM1 N_SOUT2_XI2/XI2/XI3/MM1_d N_XI2/XI2/NET17_XI2/XI2/XI3/MM1_g
+ N_VDD_XI2/XI2/XI3/MM1_s N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI2/XI0/XI2/MM1 N_XI2/XI0/NET20_XI2/XI0/XI2/MM1_d N_NET4_XI2/XI0/XI2/MM1_g
+ N_VDD_XI2/XI0/XI2/MM1_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI2/XI0/XI1/MM3 N_XI2/XI0/XI1/NET25_XI2/XI0/XI1/MM3_d
+ N_XI2/XI0/NET19_XI2/XI0/XI1/MM3_g N_XI2/XI0/XI1/NET32_XI2/XI0/XI1/MM3_s
+ N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI2/XI0/XI1/MM2 N_XI2/XI0/XI1/NET25_XI2/XI0/XI1/MM3_d N_SOUT2_XI2/XI0/XI1/MM2_g
+ N_XI2/XI0/XI1/NET26_XI2/XI0/XI1/MM2_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI2/XI0/XI1/MM5 N_XI2/XI0/XI1/NET31_XI2/XI0/XI1/MM5_d N_SOUT2_XI2/XI0/XI1/MM5_g
+ N_XI2/XI0/XI1/NET32_XI2/XI0/XI1/MM5_s N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI2/XI0/XI1/MM4 N_XI2/XI0/XI1/NET31_XI2/XI0/XI1/MM5_d
+ N_XI2/XI0/NET19_XI2/XI0/XI1/MM4_g N_XI2/XI0/XI1/NET26_XI2/XI0/XI1/MM4_s
+ N_VDD_XI2/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI2/XI0/XI1/MM11 N_XI2/XI0/XI1/NET23_XI2/XI0/XI1/MM11_d
+ N_XI2/XI0/NET19_XI2/XI0/XI1/MM11_g N_XI2/XI0/XI1/NET28_XI2/XI0/XI1/MM11_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI2/XI0/XI1/MM10 N_XI2/XI0/XI1/NET23_XI2/XI0/XI1/MM11_d
+ N_SOUT2_XI2/XI0/XI1/MM10_g N_XI2/XI0/XI1/NET22_XI2/XI0/XI1/MM10_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI2/XI0/XI1/MM13 N_XI2/XI0/XI1/NET29_XI2/XI0/XI1/MM13_d
+ N_SOUT2_XI2/XI0/XI1/MM13_g N_XI2/XI0/XI1/NET28_XI2/XI0/XI1/MM13_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI2/XI0/XI1/MM12 N_XI2/XI0/XI1/NET29_XI2/XI0/XI1/MM13_d
+ N_XI2/XI0/NET19_XI2/XI0/XI1/MM12_g N_XI2/XI0/XI1/NET22_XI2/XI0/XI1/MM12_s
+ N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI2/XI0/XI0/MM9 XI2/XI0/XI0/NET30 N_XI2/XI0/NET19_XI2/XI0/XI0/MM9_g
+ N_VDD_XI2/XI0/XI0/MM9_s N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=5.04e-14 AS=3.78e-14 PD=1e-06 PS=9.3e-07
mXI2/XI0/XI0/MM6 N_NET3_XI2/XI0/XI0/MM6_d N_XI2/XI0/NET18_XI2/XI0/XI0/MM6_g
+ XI2/XI0/XI0/NET30 N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=3.78e-14 AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI2/XI2/MM7 XI2/XI2/NET29 N_XI2/NET20_XI2/XI2/MM7_g N_VDD_XI2/XI2/MM7_s
+ N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI2/XI2/MM6 N_XI2/XI2/NET15_XI2/XI2/MM6_d N_PHI_XI2/XI2/MM6_g XI2/XI2/NET29
+ N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
mXI2/XI2/MM5 XI2/XI2/NET28 N_XI2/XI2/NET15_XI2/XI2/MM5_g N_VDD_XI2/XI2/MM5_s
+ N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI2/XI2/MM4 N_XI2/XI2/NET17_XI2/XI2/MM4_d N_XI2/XI2/NET22_XI2/XI2/MM4_g
+ XI2/XI2/NET28 N_VDD_XI2/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14
+ AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI2/XI1/MM3 XI2/XI1/NET15 N_XI2/NET21_XI2/XI1/MM3_g N_GND_XI2/XI1/MM3_s
+ N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI1/MM2 N_XI2/NET20_XI2/XI1/MM2_d N_RST_XI2/XI1/MM2_g XI2/XI1/NET15
+ N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI2/XI0/XI0/MM4 XI2/XI0/XI0/NET29 N_XI2/XI0/NET19_XI2/XI0/XI0/MM4_g
+ N_GND_XI2/XI0/XI0/MM4_s N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI2/XI0/XI0/MM1 N_NET3_XI2/XI0/XI0/MM1_d N_XI2/XI0/NET18_XI2/XI0/XI0/MM1_g
+ XI2/XI0/XI0/NET29 N_GND_XI2/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI2/XI2/MM1 XI2/XI2/NET26 N_XI2/NET20_XI2/XI2/MM1_g N_GND_XI2/XI2/MM1_s
+ N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI2/MM8 N_XI2/XI2/NET15_XI2/XI2/MM8_d N_XI2/XI2/NET22_XI2/XI2/MM8_g
+ XI2/XI2/NET26 N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14
+ AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI2/XI2/MM2 XI2/XI2/NET023 N_XI2/XI2/NET15_XI2/XI2/MM2_g N_GND_XI2/XI2/MM2_s
+ N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI2/XI2/MM0 N_XI2/XI2/NET17_XI2/XI2/MM0_d N_PHI_XI2/XI2/MM0_g XI2/XI2/NET023
+ N_GND_XI2/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI0/XI0/MM0 N_COUT_XI3/XI0/XI0/MM0_d N_XI3/XI0/NET20_XI3/XI0/XI0/MM0_g
+ N_XI3/XI0/XI0/NET15_XI3/XI0/XI0/MM0_s N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=1.8e-07 AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI3/XI0/XI0/MM3 N_XI3/XI0/XI0/NET15_XI3/XI0/XI0/MM3_d
+ N_XI3/XI0/NET19_XI3/XI0/XI0/MM3_g N_GND_XI3/XI0/XI0/MM3_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI0/XI0/MM2 N_XI3/XI0/XI0/NET15_XI3/XI0/XI0/MM3_d
+ N_XI3/XI0/NET18_XI3/XI0/XI0/MM2_g N_GND_XI3/XI0/XI0/MM2_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI1/MM0 N_XI3/NET20_XI3/XI1/MM0_d N_XI3/NET21_XI3/XI1/MM0_g
+ N_VDD_XI3/XI1/MM0_s N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI3/XI1/MM1 N_XI3/NET20_XI3/XI1/MM0_d N_RST_XI3/XI1/MM1_g N_VDD_XI3/XI1/MM1_s
+ N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI0/XI0/MM5 N_COUT_XI3/XI0/XI0/MM5_d N_XI3/XI0/NET20_XI3/XI0/XI0/MM5_g
+ N_XI3/XI0/XI0/NET17_XI3/XI0/XI0/MM5_s N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08
+ W=3.6e-07 AD=3.78e-14 AS=3.78e-14 PD=9.3e-07 PS=9.3e-07
mXI3/XI0/XI0/MM8 N_XI3/XI0/XI0/NET17_XI3/XI0/XI0/MM8_d
+ N_XI3/XI0/NET19_XI3/XI0/XI0/MM8_g N_VDD_XI3/XI0/XI0/MM8_s
+ N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI3/XI0/XI0/MM7 N_XI3/XI0/XI0/NET17_XI3/XI0/XI0/MM8_d
+ N_XI3/XI0/NET18_XI3/XI0/XI0/MM7_g N_VDD_XI3/XI0/XI0/MM7_s
+ N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI3/XI0/XI1/MM6 N_XI3/XI0/XI1/NET26_XI3/XI0/XI1/MM6_d N_A3_XI3/XI0/XI1/MM6_g
+ N_VDD_XI3/XI0/XI1/MM6_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07
+ AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI3/XI0/XI1/MM7 N_XI3/XI0/XI1/NET32_XI3/XI0/XI1/MM7_d
+ N_XI3/XI0/NET18_XI3/XI0/XI1/MM7_g N_VDD_XI3/XI0/XI1/MM7_s
+ N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=5.67e-14 AS=5.67e-14
+ PD=1.29e-06 PS=1.29e-06
mXI3/XI0/XI1/MM0 N_XI3/NET21_XI3/XI0/XI1/MM0_d N_XI3/XI0/NET20_XI3/XI0/XI1/MM0_g
+ N_XI3/XI0/XI1/NET25_XI3/XI0/XI1/MM0_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI3/XI0/XI1/MM1 N_XI3/NET21_XI3/XI0/XI1/MM1_d N_NET3_XI3/XI0/XI1/MM1_g
+ N_XI3/XI0/XI1/NET31_XI3/XI0/XI1/MM1_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=5.67e-14 AS=5.67e-14 PD=1.29e-06 PS=1.29e-06
mXI3/XI0/XI1/MM14 N_XI3/XI0/XI1/NET22_XI3/XI0/XI1/MM14_d N_A3_XI3/XI0/XI1/MM14_g
+ N_GND_XI3/XI0/XI1/MM14_s N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07
+ AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI3/XI0/XI1/MM15 N_XI3/XI0/XI1/NET28_XI3/XI0/XI1/MM15_d
+ N_XI3/XI0/NET18_XI3/XI0/XI1/MM15_g N_GND_XI3/XI0/XI1/MM15_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14
+ PD=7.5e-07 PS=7.5e-07
mXI3/XI0/XI1/MM8 N_XI3/NET21_XI3/XI0/XI1/MM8_d N_XI3/XI0/NET20_XI3/XI0/XI1/MM8_g
+ N_XI3/XI0/XI1/NET23_XI3/XI0/XI1/MM8_s N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI3/XI0/XI1/MM9 N_XI3/NET21_XI3/XI0/XI1/MM9_d N_NET3_XI3/XI0/XI1/MM9_g
+ N_XI3/XI0/XI1/NET29_XI3/XI0/XI1/MM9_s N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL
+ L=5e-08 W=2.7e-07 AD=2.835e-14 AS=2.835e-14 PD=7.5e-07 PS=7.5e-07
mXI3/XI0/XI3/MM0 N_XI3/XI0/NET18_XI3/XI0/XI3/MM0_d N_A3_XI3/XI0/XI3/MM0_g
+ N_GND_XI3/XI0/XI3/MM0_s N_GND_XI3/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI3/XI2/XI4/MM0 N_XI3/XI2/NET22_XI3/XI2/XI4/MM0_d N_PHI_XI3/XI2/XI4/MM0_g
+ N_GND_XI3/XI2/XI4/MM0_s N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI3/XI0/XI4/MM0 N_XI3/XI0/NET19_XI3/XI0/XI4/MM0_d N_SOUT3_XI3/XI0/XI4/MM0_g
+ N_GND_XI3/XI0/XI4/MM0_s N_GND_XI3/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI3/XI2/XI3/MM0 N_SOUT3_XI3/XI2/XI3/MM0_d N_XI3/XI2/NET17_XI3/XI2/XI3/MM0_g
+ N_GND_XI3/XI2/XI3/MM0_s N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI3/XI0/XI2/MM0 N_XI3/XI0/NET20_XI3/XI0/XI2/MM0_d N_NET3_XI3/XI0/XI2/MM0_g
+ N_GND_XI3/XI0/XI2/MM0_s N_GND_XI3/XI0/XI3/MM0_b NMOS_VTL L=5e-08 W=9e-08
+ AD=9.45e-15 AS=9.45e-15 PD=3.9e-07 PS=3.9e-07
mXI3/XI0/XI3/MM1 N_XI3/XI0/NET18_XI3/XI0/XI3/MM1_d N_A3_XI3/XI0/XI3/MM1_g
+ N_VDD_XI3/XI0/XI3/MM1_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI3/XI2/XI4/MM1 N_XI3/XI2/NET22_XI3/XI2/XI4/MM1_d N_PHI_XI3/XI2/XI4/MM1_g
+ N_VDD_XI3/XI2/XI4/MM1_s N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI3/XI0/XI4/MM1 N_XI3/XI0/NET19_XI3/XI0/XI4/MM1_d N_SOUT3_XI3/XI0/XI4/MM1_g
+ N_VDD_XI3/XI0/XI4/MM1_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI3/XI2/XI3/MM1 N_SOUT3_XI3/XI2/XI3/MM1_d N_XI3/XI2/NET17_XI3/XI2/XI3/MM1_g
+ N_VDD_XI3/XI2/XI3/MM1_s N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI3/XI0/XI2/MM1 N_XI3/XI0/NET20_XI3/XI0/XI2/MM1_d N_NET3_XI3/XI0/XI2/MM1_g
+ N_VDD_XI3/XI0/XI2/MM1_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=1.89e-14 PD=5.7e-07 PS=5.7e-07
mXI3/XI0/XI1/MM3 N_XI3/XI0/XI1/NET25_XI3/XI0/XI1/MM3_d
+ N_XI3/XI0/NET19_XI3/XI0/XI1/MM3_g N_XI3/XI0/XI1/NET32_XI3/XI0/XI1/MM3_s
+ N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI3/XI0/XI1/MM2 N_XI3/XI0/XI1/NET25_XI3/XI0/XI1/MM3_d N_SOUT3_XI3/XI0/XI1/MM2_g
+ N_XI3/XI0/XI1/NET26_XI3/XI0/XI1/MM2_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI3/XI0/XI1/MM5 N_XI3/XI0/XI1/NET31_XI3/XI0/XI1/MM5_d N_SOUT3_XI3/XI0/XI1/MM5_g
+ N_XI3/XI0/XI1/NET32_XI3/XI0/XI1/MM5_s N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08
+ W=5.4e-07 AD=7.56e-14 AS=5.67e-14 PD=1.36e-06 PS=1.29e-06
mXI3/XI0/XI1/MM4 N_XI3/XI0/XI1/NET31_XI3/XI0/XI1/MM5_d
+ N_XI3/XI0/NET19_XI3/XI0/XI1/MM4_g N_XI3/XI0/XI1/NET26_XI3/XI0/XI1/MM4_s
+ N_VDD_XI3/XI0/XI1/MM6_b PMOS_VTL L=5e-08 W=5.4e-07 AD=7.56e-14 AS=5.67e-14
+ PD=1.36e-06 PS=1.29e-06
mXI3/XI0/XI1/MM11 N_XI3/XI0/XI1/NET23_XI3/XI0/XI1/MM11_d
+ N_XI3/XI0/NET19_XI3/XI0/XI1/MM11_g N_XI3/XI0/XI1/NET28_XI3/XI0/XI1/MM11_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI3/XI0/XI1/MM10 N_XI3/XI0/XI1/NET23_XI3/XI0/XI1/MM11_d
+ N_SOUT3_XI3/XI0/XI1/MM10_g N_XI3/XI0/XI1/NET22_XI3/XI0/XI1/MM10_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI3/XI0/XI1/MM13 N_XI3/XI0/XI1/NET29_XI3/XI0/XI1/MM13_d
+ N_SOUT3_XI3/XI0/XI1/MM13_g N_XI3/XI0/XI1/NET28_XI3/XI0/XI1/MM13_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI3/XI0/XI1/MM12 N_XI3/XI0/XI1/NET29_XI3/XI0/XI1/MM13_d
+ N_XI3/XI0/NET19_XI3/XI0/XI1/MM12_g N_XI3/XI0/XI1/NET22_XI3/XI0/XI1/MM12_s
+ N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=2.7e-07 AD=3.78e-14 AS=2.835e-14
+ PD=8.2e-07 PS=7.5e-07
mXI3/XI0/XI0/MM9 XI3/XI0/XI0/NET30 N_XI3/XI0/NET19_XI3/XI0/XI0/MM9_g
+ N_VDD_XI3/XI0/XI0/MM9_s N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=5.04e-14 AS=3.78e-14 PD=1e-06 PS=9.3e-07
mXI3/XI0/XI0/MM6 N_COUT_XI3/XI0/XI0/MM6_d N_XI3/XI0/NET18_XI3/XI0/XI0/MM6_g
+ XI3/XI0/XI0/NET30 N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07
+ AD=3.78e-14 AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI3/XI2/MM7 XI3/XI2/NET29 N_XI3/NET20_XI3/XI2/MM7_g N_VDD_XI3/XI2/MM7_s
+ N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI3/XI2/MM6 N_XI3/XI2/NET15_XI3/XI2/MM6_d N_PHI_XI3/XI2/MM6_g XI3/XI2/NET29
+ N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14 AS=5.04e-14
+ PD=9.3e-07 PS=1e-06
mXI3/XI2/MM5 XI3/XI2/NET28 N_XI3/XI2/NET15_XI3/XI2/MM5_g N_VDD_XI3/XI2/MM5_s
+ N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=5.04e-14 AS=3.78e-14
+ PD=1e-06 PS=9.3e-07
mXI3/XI2/MM4 N_XI3/XI2/NET17_XI3/XI2/MM4_d N_XI3/XI2/NET22_XI3/XI2/MM4_g
+ XI3/XI2/NET28 N_VDD_XI3/XI2/XI4/MM1_b PMOS_VTL L=5e-08 W=3.6e-07 AD=3.78e-14
+ AS=5.04e-14 PD=9.3e-07 PS=1e-06
mXI3/XI1/MM3 XI3/XI1/NET15 N_XI3/NET21_XI3/XI1/MM3_g N_GND_XI3/XI1/MM3_s
+ N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI1/MM2 N_XI3/NET20_XI3/XI1/MM2_d N_RST_XI3/XI1/MM2_g XI3/XI1/NET15
+ N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
mXI3/XI0/XI0/MM4 XI3/XI0/XI0/NET29 N_XI3/XI0/NET19_XI3/XI0/XI0/MM4_g
+ N_GND_XI3/XI0/XI0/MM4_s N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=2.52e-14 AS=1.89e-14 PD=6.4e-07 PS=5.7e-07
mXI3/XI0/XI0/MM1 N_COUT_XI3/XI0/XI0/MM1_d N_XI3/XI0/NET18_XI3/XI0/XI0/MM1_g
+ XI3/XI0/XI0/NET29 N_GND_XI3/XI0/XI1/MM14_b NMOS_VTL L=5e-08 W=1.8e-07
+ AD=1.89e-14 AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI3/XI2/MM1 XI3/XI2/NET26 N_XI3/NET20_XI3/XI2/MM1_g N_GND_XI3/XI2/MM1_s
+ N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI2/MM8 N_XI3/XI2/NET15_XI3/XI2/MM8_d N_XI3/XI2/NET22_XI3/XI2/MM8_g
+ XI3/XI2/NET26 N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14
+ AS=2.52e-14 PD=5.7e-07 PS=6.4e-07
mXI3/XI2/MM2 XI3/XI2/NET023 N_XI3/XI2/NET15_XI3/XI2/MM2_g N_GND_XI3/XI2/MM2_s
+ N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=2.52e-14 AS=1.89e-14
+ PD=6.4e-07 PS=5.7e-07
mXI3/XI2/MM0 N_XI3/XI2/NET17_XI3/XI2/MM0_d N_PHI_XI3/XI2/MM0_g XI3/XI2/NET023
+ N_GND_XI3/XI2/XI4/MM0_b NMOS_VTL L=5e-08 W=1.8e-07 AD=1.89e-14 AS=2.52e-14
+ PD=5.7e-07 PS=6.4e-07
*
.include "4_bit_accumulator.pex.netlist.4_BIT_ACCUMULATOR.pxi"
*
.ends
*
*
x1 GND PHI RST VDD CIN COUT A0 SOUT0 A1 SOUT1 A2 SOUT2 A3 SOUT3 four_bit_accumulator

*------------------------------------------------------------------------
* Stimulus
*------------------------------------------------------------------------

.tran 1ps 1820ps SWEEP clk_period POI 1 100


.END